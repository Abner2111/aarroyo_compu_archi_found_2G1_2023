module PWM_tb();

	reg [3:0] Porcentaje;
	reg SLK;
	wire pwm;
	
	PWM_module test(.Porcentaje(Porcentaje), .SLK(SLK), .pwm(pwm));
	
	initial begin
	
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
		#1 SLK = ~SLK;
	
	end
	
	initial begin

		SLK = 0;
		Porcentaje = 1;
		#10
		Porcentaje = 2;
		#10
		Porcentaje = 3;
		#10;
		Porcentaje = 4;
		#10;
		Porcentaje = 5;
		#10;
		Porcentaje = 6;
		#10;
		Porcentaje = 7;
		#10;
		Porcentaje = 8;
		#10;
		Porcentaje = 9;
		#10;
		Porcentaje = 10;
		#10;
		Porcentaje = 0;
		#10;
		Porcentaje = 1;
		#10
		Porcentaje = 2;
		#10
		Porcentaje = 3;
		#10;
		Porcentaje = 4;
		#10;
		Porcentaje = 5;
		#10;
		Porcentaje = 6;
		#10;
		Porcentaje = 7;
		#10;
		Porcentaje = 8;
		#10;
		Porcentaje = 9;
		#10;
		Porcentaje = 10;
		#10;
	
	$finish; // Termina la simulación
	end

endmodule